------------------------------
-- Elementos de Sistemas
-- Avaliacao Pratica 1
--
-- 10/2019
--
-- Questão 5
------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity questao2 is
  port (
    a  : in  STD_LOGIC_VECTOR(7 downto 0);
    sel: in  STD_LOGIC_VECTOR(1 downto 0);
    b  : out STD_LOGIC_VECTOR(3 downto 0));
end entity;

architecture  rtl OF questao2 IS

begin

end architecture;
